library IEEE;
use IEEE.std_logic_1164.all;

entity tb_N_bitRegister is
  generic(gCLK_HPER   : time := 50 ns;
		N			: integer := 32);
end tb_N_bitRegister;

architecture behavior of tb_N_bitRegister is
  
  constant cCLK_PER  : time := gCLK_HPER * 2;

  component N_bitRegister
    port(i_CLK        : in std_logic;     		-- Clock input
         i_RST        : in std_logic;     		-- Reset input
         i_WE         : in std_logic;     		-- Write enable input
         i_D          : in std_logic_vector(N-1 downto 0);     -- Data value input
         o_Q          : out std_logic_vector(N-1 downto 0));   -- Data value output
  end component;


  signal s_CLK, s_RST, s_WE  : std_logic;
  signal s_D, s_Q : std_logic_vector(N-1 downto 0);

begin

  DUT: N_bitRegister
  port map(i_CLK => s_CLK, 
           i_RST => s_RST,
           i_WE  => s_WE,
           i_D   => s_D,
           o_Q   => s_Q);

  P_CLK: process
  begin
    s_CLK <= '0';
    wait for gCLK_HPER;
    s_CLK <= '1';
    wait for gCLK_HPER;
  end process;
  
 
  P_TB: process
  begin

    s_RST <= '1';
    s_WE  <= '0';
    s_D   <= "00000000000000000000000000000000";
    wait for cCLK_PER;

    s_RST <= '0';
    s_WE  <= '1';
    s_D   <= "11111111111111111111111111111111";
    wait for cCLK_PER;  

    s_RST <= '0';
    s_WE  <= '0';
    s_D   <= "00000000000000000000000000000000";
    wait for cCLK_PER;  


    s_RST <= '0';
    s_WE  <= '1';
    s_D   <= "00000000000000000000000000000011";
    wait for cCLK_PER;  


    s_RST <= '0';
    s_WE  <= '0';
    s_D   <= "11111111111111111111111111111111";
    wait for cCLK_PER;  
	

    s_RST <= '1';
    s_WE  <= '0';
    s_D   <= "11111111111111111111111111111111";
    wait for cCLK_PER;

    wait;
  end process;
  
end behavior;