library IEEE;
use IEEE.std_logic_1164.all;

use work.mypack.all;

entity tb_mux32t1 is
  generic(gCLK_HPER : time := 50 ns);  
end tb_mux32t1;

architecture behavior of tb_mux32t1 is 
  constant cCLK_PER : time := gCLK_HPER * 2;

  component mux32t1
    port(
      i_I : in TwoDArray;                     -- 32 inputs
      i_S : in std_logic_vector(4 downto 0);  -- Select input (5-bit)
      o_O : out std_logic_vector(31 downto 0) -- Output (32-bit)
    );
  end component;

  -- Signal declarations for connecting to the multiplexer
  signal s_I : TwoDArray;
  signal s_S : std_logic_vector(4 downto 0);
  signal s_O : std_logic_vector(31 downto 0);

begin
  -- Instantiate the multiplexer component
  DUT: mux32t1
    port map(i_I => s_I, i_S => s_S, o_O => s_O);

  -- Initialization process to set input data
  P_INIT: process
  begin
    -- Initialize all inputs to 0
    for i in 0 to 31 loop
      s_I(i) <= (others => '0');
    end loop;
    wait for cCLK_PER * 4;

    -- Set different values for testing
    for i in 10 to 20 loop
      s_I(i) <= (others => '1');  -- Inputs 10-20 set to all 1's
    end loop;
    for i in 20 to 31 loop
      s_I(i) <= (others => '1');  -- Inputs 21-31 set to all 1's
    end loop;

    wait;
  end process;

  -- Testbench process to apply test vectors
  P_TB: process
  begin
    -- Test Case 1 --
    s_S <= "00001";
    wait for cCLK_PER; 
	
    -- Test Case 2 --
    s_S <= "00100";
    wait for cCLK_PER; 
	
    -- Test Case 3 --
    s_S <= "01011";
    wait for cCLK_PER; 
	
    -- Test Case 4 --
    s_S <= "11111";
    wait for cCLK_PER;

    wait;
  end process;
end behavior;
