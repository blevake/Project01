library IEEE;
use IEEE.std_logic_1164.all;

entity tb_regfile is
  generic(gCLK_HPER : time := 50 ns);  
end tb_regfile;

architecture behavior of tb_regfile is
  constant cCLK_PER : time := gCLK_HPER * 2;

  component regfile
    port(
      clk    : in std_logic;
      i_wA   : in std_logic_vector(4 downto 0);  -- Write address
      i_rA0  : in std_logic_vector(4 downto 0);  -- Read address 0
      i_rA1  : in std_logic_vector(4 downto 0);  -- Read address 1
      i_wD   : in std_logic_vector(31 downto 0); -- Write data
      i_wE   : in std_logic;                     -- Write enable
      o_RD0  : out std_logic_vector(31 downto 0);-- Read data 0
      o_RD1  : out std_logic_vector(31 downto 0) -- Read data 1
    );
  end component;

  -- Signals for connecting to the register file
  signal s_CLK : std_logic;
  signal s_wA, s_rA0, s_rA1 : std_logic_vector(4 downto 0);
  signal s_wD, s_oRD0, s_oRD1 : std_logic_vector(31 downto 0);
  signal s_wE : std_logic;

begin
  -- Instantiate the register file component
  DUT: regfile
    port map(
      clk   => s_CLK,
      i_wA  => s_wA,
      i_rA0 => s_rA0,
      i_rA1 => s_rA1,
      i_wD  => s_wD,
      i_wE  => s_wE,
      o_RD0 => s_oRD0,
      o_RD1 => s_oRD1
    );

  -- Clock generation process
  P_CLK: process
  begin
    s_CLK <= '0';
    wait for gCLK_HPER;
    s_CLK <= '1';
    wait for gCLK_HPER;
  end process;
  
  P_TB: process
  begin
    -- Test Case 1 --
    s_wA <= "00001";  -- Write address = 1
    s_rA0 <= "00001"; -- Read address 0 = 1
    s_rA1 <= "00010"; -- Read address 1 = 2
    s_wD <= x"00000003";  -- Write data = 3
    s_wE <= '1';          -- Write enable
    wait for cCLK_PER;  -- Expected Output: Register 1 = 3, others = 0

    -- Test Case 2 --
    s_wE <= '0';          -- Disable write
    wait for cCLK_PER;    -- Expected Output: Register 1 = 3, others = 0

    -- Test Case 3 --
    s_wA <= "00010";      -- Write address = 2
    s_wD <= x"0000000F";  -- Write data = 15
    s_wE <= '1';          -- Write enable
    wait for cCLK_PER;    -- Expected Output: Register 2 = 15, register 1 = 3

    -- Test Case 4 --
    s_wE <= '0';          -- Disable write
    wait for cCLK_PER;    -- Expected Output: Registers hold values

    wait;
  end process;
end behavior;
